`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Mohammad Musawer
// 
// Create Date: 08/05/2021 02:40:10 PM
// Project Name: Central Processing Unit Design in Verilog
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module control_unit(

    );
endmodule


module ALU(

    );
endmodule


module RAM(

    );
endmodule


module register(

    );
endmodule
